`ifndef INTERFACE_SV
`define INTERFACE_SV
interface intf;
  logic [2:0]in;
  logic [7:0]out;
endinterface
`endif